library verilog;
use verilog.vl_types.all;
entity Pipline is
end Pipline;
