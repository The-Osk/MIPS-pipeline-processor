library verilog;
use verilog.vl_types.all;
entity ALU_Test is
end ALU_Test;
