library verilog;
use verilog.vl_types.all;
entity CLK is
    port(
        clk             : out    vl_logic
    );
end CLK;
