library verilog;
use verilog.vl_types.all;
entity Test_Reg_File is
end Test_Reg_File;
