library verilog;
use verilog.vl_types.all;
entity Top_Module is
    port(
        x               : in     vl_logic;
        y               : out    vl_logic
    );
end Top_Module;
