library verilog;
use verilog.vl_types.all;
entity Pipline2 is
    port(
        initial_PC      : in     vl_logic_vector(31 downto 0)
    );
end Pipline2;
