library verilog;
use verilog.vl_types.all;
entity Test_CLK is
end Test_CLK;
