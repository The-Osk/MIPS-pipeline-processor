module Top_Module(x,y);
/*
reg [31:0]initial_PC;
Pipline2 Pipline21(initial_PC);
initial
begin
initial_PC=0;
#1 $display("hahha = %h",Pipline21.Reg_File1);
end

*/
input x;
output y;
endmodule
