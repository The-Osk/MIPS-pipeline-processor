library verilog;
use verilog.vl_types.all;
entity Test_Data_Mem is
end Test_Data_Mem;
