library verilog;
use verilog.vl_types.all;
entity Test_PC_Add4 is
end Test_PC_Add4;
