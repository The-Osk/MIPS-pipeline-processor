library verilog;
use verilog.vl_types.all;
entity Test_Instruc_mem is
end Test_Instruc_mem;
